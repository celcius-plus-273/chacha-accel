module serializer
#(

)
(

);

endmodule