/**
 *  ARX operation implementation
 */