module chacha_accel (

)


endmodule